

module maquina_cafe(input clk, rst, e, l, x, m, a, C, Q,
						  output bebidaLista, agua, cafe, leche, choco, azucar,
						  output [6:0] hex1, hex2);
						  
endmodule 